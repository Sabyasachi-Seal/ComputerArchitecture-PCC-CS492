----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:06:10 06/14/2022 
-- Design Name: 
-- Module Name:    xor_rtl - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity xor_rtl is
    Port ( xa : in  STD_LOGIC;
           xb : in  STD_LOGIC;
           xout : out  STD_LOGIC);
end xor_rtl;

architecture Behavioral of xor_rtl is

begin
xout <= ((not xa) and xb) or ((not xb) and xa);

end Behavioral;

